// EXECUTE CYCLE CODE:
//module execute cycle-------------------------------------------------------------------
module execute_cycle(clk, rst, RegWriteE, ALUSrcE, MemWriteE, ResultSrcE, BranchE, ALUControlE, RD1_E, RD2_E, Imm_Ext_E, RD_E, PCE, PCPlus4E, PCTargetE, PCSrcE, RegWriteM, MemWriteM, ResultSrcM, RD_M, PCPlus4M, WriteDataM, ALUResultM);

input clk, rst;
input RegWriteE, ALUSrcE, MemWriteE, ResultSrcE, BranchE;
input [2:0] ALUControlE;
input [31:0] RD1_E, RD2_E, Imm_Ext_E;
input [4:0] RD_E;
input [31:0] PCE, PCPlus4E;
output [31:0] PCTargetE, ALUResultM, WriteDataM, PCPlus4M;
output PCSrcE, RegWriteM, MemWriteM, ResultSrcM;
output[4:0] RD_M;

//declare interim wires:
wire [31:0] Src_b, Result_E;
wire zero_E;

//declaration of modules:
ALU alu(.A(RD1_E),
        .B(Src_b),
        .Result(Result_E),
        .ALUControl(ALUControlE),
        .OverFlow(),
        .Carry(),
        .Zero(zero_E),
        .Negative());

Mux alu_src_mux(.a(RD2_E),
                .b(Imm_Ext_E), 
                .s(ALUSrcE),
                .c(Src_b));

PC_Adder branch_adder(.a(PCE),
                      .b(Imm_Ext_E),
                      .c(PCTargetE));

//declaration of registers:
reg RegWriteE_r, MemWriteE_r, ResultSrcE_r;
reg [4:0] RD_E_r;
reg [31:0] PCPlus4E_r, RD2_E_r, ResultE_r;

always @(posedge clk or posedge rst) begin 
if(rst==1'b1) begin 
    RegWriteE_r<=1'b0;
    MemWriteE_r<=1'b0;
    ResultSrcE_r<=1'b0;
    RD_E_r<=5'b0;
    PCPlus4E_r<=32'b0;
    RD2_E_r<=32'b0;
    ResultE_r<=32'b0;
   end
else begin 
    RegWriteE_r<=RegWriteE;
    MemWriteE_r<=MemWriteE;
    ResultSrcE_r<=ResultSrcE;
    RD_E_r<=RD_E;
    PCPlus4E_r<=PCPlus4E;
    RD2_E_r<=RD2_E;
    ResultE_r<=Result_E;     
    end
end

//output assignments;
assign PCSrcE=zero_E & BranchE;
assign RegWriteM=RegWriteE_r;
assign MemWriteM=MemWriteE_r;
assign ResultSrcM=ResultSrcE_r;
assign RD_M=RD_E_r;
assign PCPlus4M=PCPlus4E_r;
assign WriteDataM=RD2_E_r;
assign ALUResultM=ResultE_r;
endmodule
